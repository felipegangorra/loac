// Felipe Gangorra - UFCG
// Meu primeiro código em SystemVeriLog

module HelloWorld();
  initial begin
    $display("Hello, World!");
  end
endmodule